library verilog;
use verilog.vl_types.all;
entity zero_testbench is
end zero_testbench;
